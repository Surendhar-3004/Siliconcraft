interface inter;
  logic clk;
 // logic reset;
  logic [3:0]wdata;
  logic [3:0]addr;
  logic w_en;
  logic [3:0]rdata;
  
endinterface
