module NAND_gate(output Y, input A, B);
  nand(Y, A, B);
endmodule;
