interface inter;
  logic a;
  logic b;
  logic cin;
  logic sum;
  logic cout;
endinterface
