class transaction;
  
  bit clk;
  bit rst;
  rand logic d;
  reg q;
  //constraint cs{ inside [d!=d;]}
endclass
