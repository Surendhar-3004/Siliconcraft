class transaction;
  rand bit a;
  rand bit b;
  rand bit cin;
  bit sum;
  bit cout;
endclass
