module nor_gate(output Y, input A, B);
  nor(Y, A, B);
endmodule;
