module AND_gate(output Y, input A, B);
  and(Y, A, B);
endmodule
