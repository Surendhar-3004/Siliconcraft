module not_gate(
  input a,
  output b);
  not(b,a);
endmodule
