module xnor_gate(
  input A,
  input B,
  output Y);
  xnor(Y,A,B);
endmodule
