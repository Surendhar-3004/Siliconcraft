class transaction;
  bit clk;
 // bit reset;
  rand bit [3:0]wdata;
  rand bit [3:0]addr;
  bit w_en;
  reg rdata;
endclass
